// and2.v  M.L. Johnston
// 2-Input AND Gate

module and2(	input a,b,
		output y);
	
	assign y = a & b;
	
endmodule

