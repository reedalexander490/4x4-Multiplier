// or2.v  Hugo Korte
// 2-Input or Gate

module or2(	input a,b,
		output y);
	
	assign y = a | b;
	
endmodule

